module Qb(D, clk, O);
endmodule
